module encoder_10to4_tb;

    reg  [9:0] d;
    wire [3:0] y;

    encoder_10to4 dut(.d(d), .y(y));

    initial begin

        d = 10'b0000000001; #10;
        d = 10'b0000000010; #10;
        d = 10'b0000000100; #10;
        d = 10'b0000001000; #10;
        d = 10'b0000010000; #10;
        d = 10'b0000100000; #10;
        d = 10'b0001000000; #10;
        d = 10'b0010000000; #10;
        d = 10'b0100000000; #10;
        d = 10'b1000000000; #10;

        $finish;
    end

endmodule
