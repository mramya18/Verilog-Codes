module ripple_carry_adder_tb;
reg [3:0]a,b;
reg cin;
wire [2:0]s;
wire cout;

ripple_carry_adder dut(.a(a), .b(b), .cin(cin), .s(s), .cout(cout));
initial begin
a=4'b0000; b= 4'b0000; cin=0; #10;
a=4'b0001; b= 4'b0001; cin=0; #10;
a=4'b0010; b= 4'b0010; cin=0; #10;
a=4'b0011; b= 4'b0011; cin=0; #10;
a=4'b0100; b= 4'b0100; cin=0; #10;
a=4'b0101; b= 4'b0101; cin=0; #10;
a=4'b0110; b= 4'b0110; cin=0; #10;
a=4'b0111; b= 4'b0111; cin=0; #10;
a=4'b1000; b= 4'b1000; cin=0; #10;
a=4'b1001; b= 4'b1001; cin=0; #10;
a=4'b1010; b= 4'b1010; cin=0; #10;
a=4'b1011; b= 4'b1011; cin=0; #10;
a=4'b1100; b= 4'b1100; cin=0; #10;
a=4'b1101; b= 4'b1101; cin=0; #10;
a=4'b1110; b= 4'b1110; cin=0; #10;
a=4'b1111; b= 4'b1111; cin=0; #10;

$finish;
end


endmodule
